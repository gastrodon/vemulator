module main

const (
	nop    = 0x00
	lxi_b  = 0x01
	stax_b = 0x02
	inx_b  = 0x03
	inr_b  = 0x04
	dcr_b  = 0x05
	mvi_b  = 0x06
	rcl    = 0x07
	dad_b  = 0x09
	sta    = 0x32
	lda    = 0x3a
	inr_a  = 0x3c
)
